 // ---------- SEQUENCER -----------------
  typedef uvm_sequencer #(my_txn) my_sqr ;
